package seq_pkg;

    import uvm_pkg::*;
    import ahb_pkg::*;

    `include "ahb_read_sequence.sv"
    `include "ahb_write_sequence.sv"

endpackage